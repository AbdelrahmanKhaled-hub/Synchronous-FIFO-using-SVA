package FIFO_shared_pkg;

int Error_count=0,Correct_count=0;
bit test_finished=0;

endpackage
